-- pll25.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pll25 is
	port (
		ref_clk_clk        : in  std_logic := '0'; --      ref_clk.clk
		ref_reset_reset    : in  std_logic := '0'; --    ref_reset.reset
		reset_source_reset : out std_logic;        -- reset_source.reset
		vga_clk_clk        : out std_logic         --      vga_clk.clk
	);
end entity pll25;

architecture rtl of pll25 is
	component pll25_video_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			vga_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component pll25_video_pll_0;

begin

	video_pll_0 : component pll25_video_pll_0
		port map (
			ref_clk_clk        => ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => ref_reset_reset,    --    ref_reset.reset
			vga_clk_clk        => vga_clk_clk,        --      vga_clk.clk
			reset_source_reset => reset_source_reset  -- reset_source.reset
		);

end architecture rtl; -- of pll25
